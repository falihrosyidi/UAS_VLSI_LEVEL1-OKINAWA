`ifndef TANH
`define TANH

module tanh #(
    parameter WIDTH = 32
) (
    input [WIDTH-1:0] a,
    output [WIDTH-1:0] y
);
    // algoritma tanh
endmodule

`endif 