`ifndef SIGMOID
`define SIGMOID

module sigmoid #(
    parameter WIDTH = 32
) (
    input [WIDTH-1:0] a,
    output [WIDTH-1:0] y
);
    // algoritma SIGMOID
endmodule

`endif 